//////////////////////////////////////////////////////////////////////////////////
//
// This file is part of the N64 RGB/YPbPr DAC project.
//
// Copyright (C) 2015-2024 by Peter Bartmann <borti4938@gmail.com>
//
// N64 RGB/YPbPr DAC is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <http://www.gnu.org/licenses/>.
//
//////////////////////////////////////////////////////////////////////////////////
//
// Company: Circuit-Board.de
// Engineer: borti4938
//
// VH-file Name:   n64adv2_hw_cfg.vh
// Project Name:   N64 Advanced Mod
// Target Devices: several devices
// Tool versions:  Altera Quartus Prime
// Description:
//
//////////////////////////////////////////////////////////////////////////////////


`ifndef _n64adv2_hw_cfg_vh_
`define _n64adv2_hw_cfg_vh_

  parameter [3:0] hdl_fw_main = 4'd2;
  parameter [7:0] hdl_fw_sub  = 8'd15;
  
//  parameter osd_font_rom_version = "V1";
  parameter osd_font_rom_version = "V2";
  parameter osd_window_color = "Darkblue";  // allowed/implemented: White, Grey, Black, Darkblue
  
//  `define VIDEO_USE_FAST_OUTPUT_REGs

`endif