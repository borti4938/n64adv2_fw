//////////////////////////////////////////////////////////////////////////////////
//
// This file is part of the N64 RGB/YPbPr DAC project.
//
// Copyright (C) 2015-2023 by Peter Bartmann <borti4938@gmail.com>
//
// N64 RGB/YPbPr DAC is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <http://www.gnu.org/licenses/>.
//
//////////////////////////////////////////////////////////////////////////////////
//
// Company:  Circuit-Board.de
// Engineer: borti4938
//
// Module Name:    font_rom_v2
// Project Name:   N64 Advanced RGB/YPbPr DAC Mod
// Target Devices: Max10, Cyclone IV and Cyclone 10 LP devices
// Tool versions:  Altera Quartus Prime
// Description:    simple line-multiplying
//
// Features: ip independent implementation of font rom
//
// This file is auto generated by script/font2rom.m
//
//////////////////////////////////////////////////////////////////////////////////


module font_rom_v2(
  CLK,
  nRST,
  char_addr,
  char_line,
  rden,
  rddata
);

input       CLK;
input       nRST;
input [6:0] char_addr;
input [3:0] char_line;
input       rden;

output reg [7:0] rddata = 8'h0;


reg [7:0] rddata_opt [0:3];
initial begin
  rddata_opt[0] = 8'h0;
  rddata_opt[1] = 8'h0;
  rddata_opt[2] = 8'h0;
  rddata_opt[3] = 8'h0;
end
reg [1:0] lsb_addr_r = 2'h00;
reg           rden_r = 1'b0;

always @(posedge CLK or negedge nRST)
  if (!nRST) begin
    rddata <= 8'h0;
    rddata_opt[0] = 8'h0;
    rddata_opt[1] = 8'h0;
    rddata_opt[2] = 8'h0;
    rddata_opt[3] = 8'h0;
    lsb_addr_r <= 2'h00;
    rden_r <= 1'b0;
  end else begin
    lsb_addr_r <= char_addr[1:0];
    rden_r <= rden;
  
    if (rden) begin
      case ({char_line,char_addr[6:2]})
        0023: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 008;
            rddata_opt[3] <= 000;
          end
        0024: begin
            rddata_opt[0] <= 012;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0034: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 028;
            rddata_opt[3] <= 000;
          end
        0036: begin
            rddata_opt[0] <= 064;
            rddata_opt[1] <= 001;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0040: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0042: begin
            rddata_opt[0] <= 048;
            rddata_opt[1] <= 006;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0044: begin
            rddata_opt[0] <= 062;
            rddata_opt[1] <= 008;
            rddata_opt[2] <= 030;
            rddata_opt[3] <= 030;
          end
        0045: begin
            rddata_opt[0] <= 048;
            rddata_opt[1] <= 063;
            rddata_opt[2] <= 028;
            rddata_opt[3] <= 127;
          end
        0046: begin
            rddata_opt[0] <= 030;
            rddata_opt[1] <= 030;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0047: begin
            rddata_opt[0] <= 048;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 006;
            rddata_opt[3] <= 030;
          end
        0048: begin
            rddata_opt[0] <= 062;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 063;
            rddata_opt[3] <= 060;
          end
        0049: begin
            rddata_opt[0] <= 031;
            rddata_opt[1] <= 127;
            rddata_opt[2] <= 127;
            rddata_opt[3] <= 060;
          end
        0050: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 030;
            rddata_opt[2] <= 120;
            rddata_opt[3] <= 103;
          end
        0051: begin
            rddata_opt[0] <= 015;
            rddata_opt[1] <= 099;
            rddata_opt[2] <= 099;
            rddata_opt[3] <= 028;
          end
        0052: begin
            rddata_opt[0] <= 063;
            rddata_opt[1] <= 028;
            rddata_opt[2] <= 063;
            rddata_opt[3] <= 030;
          end
        0053: begin
            rddata_opt[0] <= 063;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 099;
          end
        0054: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 127;
            rddata_opt[3] <= 060;
          end
        0055: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 060;
            rddata_opt[2] <= 028;
            rddata_opt[3] <= 000;
          end
        0056: begin
            rddata_opt[0] <= 012;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 007;
            rddata_opt[3] <= 000;
          end
        0057: begin
            rddata_opt[0] <= 056;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 028;
            rddata_opt[3] <= 000;
          end
        0058: begin
            rddata_opt[0] <= 007;
            rddata_opt[1] <= 024;
            rddata_opt[2] <= 048;
            rddata_opt[3] <= 007;
          end
        0059: begin
            rddata_opt[0] <= 030;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0066: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 034;
            rddata_opt[3] <= 000;
          end
        0068: begin
            rddata_opt[0] <= 096;
            rddata_opt[1] <= 003;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0072: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 030;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0074: begin
            rddata_opt[0] <= 024;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0075: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 064;
          end
        0076: begin
            rddata_opt[0] <= 099;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 051;
          end
        0077: begin
            rddata_opt[0] <= 056;
            rddata_opt[1] <= 003;
            rddata_opt[2] <= 006;
            rddata_opt[3] <= 099;
          end
        0078: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0079: begin
            rddata_opt[0] <= 024;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 012;
            rddata_opt[3] <= 051;
          end
        0080: begin
            rddata_opt[0] <= 099;
            rddata_opt[1] <= 030;
            rddata_opt[2] <= 102;
            rddata_opt[3] <= 102;
          end
        0081: begin
            rddata_opt[0] <= 054;
            rddata_opt[1] <= 070;
            rddata_opt[2] <= 102;
            rddata_opt[3] <= 102;
          end
        0082: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 048;
            rddata_opt[3] <= 102;
          end
        0083: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 119;
            rddata_opt[2] <= 099;
            rddata_opt[3] <= 054;
          end
        0084: begin
            rddata_opt[0] <= 102;
            rddata_opt[1] <= 054;
            rddata_opt[2] <= 102;
            rddata_opt[3] <= 051;
          end
        0085: begin
            rddata_opt[0] <= 045;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 099;
          end
        0086: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 115;
            rddata_opt[3] <= 012;
          end
        0087: begin
            rddata_opt[0] <= 001;
            rddata_opt[1] <= 048;
            rddata_opt[2] <= 054;
            rddata_opt[3] <= 000;
          end
        0088: begin
            rddata_opt[0] <= 024;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 006;
            rddata_opt[3] <= 000;
          end
        0089: begin
            rddata_opt[0] <= 048;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 054;
            rddata_opt[3] <= 000;
          end
        0090: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 024;
            rddata_opt[2] <= 048;
            rddata_opt[3] <= 006;
          end
        0091: begin
            rddata_opt[0] <= 024;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0093: begin
            rddata_opt[0] <= 004;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0098: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 093;
            rddata_opt[3] <= 000;
          end
        0099: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 099;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0100: begin
            rddata_opt[0] <= 112;
            rddata_opt[1] <= 007;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0102: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 012;
            rddata_opt[3] <= 024;
          end
        0104: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 030;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0105: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 035;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0106: begin
            rddata_opt[0] <= 012;
            rddata_opt[1] <= 024;
            rddata_opt[2] <= 102;
            rddata_opt[3] <= 024;
          end
        0107: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 096;
          end
        0108: begin
            rddata_opt[0] <= 115;
            rddata_opt[1] <= 015;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 048;
          end
        0109: begin
            rddata_opt[0] <= 060;
            rddata_opt[1] <= 003;
            rddata_opt[2] <= 003;
            rddata_opt[3] <= 099;
          end
        0110: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 028;
            rddata_opt[3] <= 028;
          end
        0111: begin
            rddata_opt[0] <= 012;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 024;
            rddata_opt[3] <= 048;
          end
        0112: begin
            rddata_opt[0] <= 099;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 102;
            rddata_opt[3] <= 099;
          end
        0113: begin
            rddata_opt[0] <= 102;
            rddata_opt[1] <= 006;
            rddata_opt[2] <= 070;
            rddata_opt[3] <= 099;
          end
        0114: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 048;
            rddata_opt[3] <= 054;
          end
        0115: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 127;
            rddata_opt[2] <= 103;
            rddata_opt[3] <= 099;
          end
        0116: begin
            rddata_opt[0] <= 102;
            rddata_opt[1] <= 099;
            rddata_opt[2] <= 102;
            rddata_opt[3] <= 051;
          end
        0117: begin
            rddata_opt[0] <= 012;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 099;
          end
        0118: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 025;
            rddata_opt[3] <= 012;
          end
        0119: begin
            rddata_opt[0] <= 003;
            rddata_opt[1] <= 048;
            rddata_opt[2] <= 099;
            rddata_opt[3] <= 000;
          end
        0120: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 006;
            rddata_opt[3] <= 000;
          end
        0121: begin
            rddata_opt[0] <= 048;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 006;
            rddata_opt[3] <= 000;
          end
        0122: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 006;
          end
        0123: begin
            rddata_opt[0] <= 024;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0125: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0130: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 069;
            rddata_opt[3] <= 000;
          end
        0131: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 054;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0132: begin
            rddata_opt[0] <= 124;
            rddata_opt[1] <= 031;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0134: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 006;
            rddata_opt[3] <= 048;
          end
        0136: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 030;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0137: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0138: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 048;
            rddata_opt[2] <= 060;
            rddata_opt[3] <= 024;
          end
        0139: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 048;
          end
        0140: begin
            rddata_opt[0] <= 123;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 048;
            rddata_opt[3] <= 048;
          end
        0141: begin
            rddata_opt[0] <= 054;
            rddata_opt[1] <= 003;
            rddata_opt[2] <= 003;
            rddata_opt[3] <= 096;
          end
        0142: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 028;
            rddata_opt[3] <= 028;
          end
        0143: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 126;
            rddata_opt[2] <= 048;
            rddata_opt[3] <= 024;
          end
        0144: begin
            rddata_opt[0] <= 123;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 102;
            rddata_opt[3] <= 003;
          end
        0145: begin
            rddata_opt[0] <= 102;
            rddata_opt[1] <= 038;
            rddata_opt[2] <= 038;
            rddata_opt[3] <= 003;
          end
        0146: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 048;
            rddata_opt[3] <= 054;
          end
        0147: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 127;
            rddata_opt[2] <= 111;
            rddata_opt[3] <= 099;
          end
        0148: begin
            rddata_opt[0] <= 102;
            rddata_opt[1] <= 099;
            rddata_opt[2] <= 102;
            rddata_opt[3] <= 003;
          end
        0149: begin
            rddata_opt[0] <= 012;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 099;
          end
        0150: begin
            rddata_opt[0] <= 030;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 024;
            rddata_opt[3] <= 012;
          end
        0151: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 048;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0152: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 030;
            rddata_opt[2] <= 062;
            rddata_opt[3] <= 030;
          end
        0153: begin
            rddata_opt[0] <= 062;
            rddata_opt[1] <= 030;
            rddata_opt[2] <= 006;
            rddata_opt[3] <= 110;
          end
        0154: begin
            rddata_opt[0] <= 054;
            rddata_opt[1] <= 030;
            rddata_opt[2] <= 060;
            rddata_opt[3] <= 102;
          end
        0155: begin
            rddata_opt[0] <= 024;
            rddata_opt[1] <= 063;
            rddata_opt[2] <= 031;
            rddata_opt[3] <= 030;
          end
        0156: begin
            rddata_opt[0] <= 059;
            rddata_opt[1] <= 110;
            rddata_opt[2] <= 055;
            rddata_opt[3] <= 030;
          end
        0157: begin
            rddata_opt[0] <= 063;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 099;
          end
        0158: begin
            rddata_opt[0] <= 099;
            rddata_opt[1] <= 102;
            rddata_opt[2] <= 063;
            rddata_opt[3] <= 000;
          end
        0162: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 069;
            rddata_opt[3] <= 000;
          end
        0163: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 028;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0164: begin
            rddata_opt[0] <= 127;
            rddata_opt[1] <= 127;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0166: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 127;
            rddata_opt[3] <= 127;
          end
        0168: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0169: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 024;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0170: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 048;
            rddata_opt[2] <= 255;
            rddata_opt[3] <= 126;
          end
        0171: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 127;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 024;
          end
        0172: begin
            rddata_opt[0] <= 107;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 024;
            rddata_opt[3] <= 028;
          end
        0173: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 031;
            rddata_opt[2] <= 031;
            rddata_opt[3] <= 048;
          end
        0174: begin
            rddata_opt[0] <= 030;
            rddata_opt[1] <= 062;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0175: begin
            rddata_opt[0] <= 003;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 096;
            rddata_opt[3] <= 012;
          end
        0176: begin
            rddata_opt[0] <= 123;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 062;
            rddata_opt[3] <= 003;
          end
        0177: begin
            rddata_opt[0] <= 102;
            rddata_opt[1] <= 062;
            rddata_opt[2] <= 062;
            rddata_opt[3] <= 003;
          end
        0178: begin
            rddata_opt[0] <= 063;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 048;
            rddata_opt[3] <= 030;
          end
        0179: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 107;
            rddata_opt[2] <= 127;
            rddata_opt[3] <= 099;
          end
        0180: begin
            rddata_opt[0] <= 062;
            rddata_opt[1] <= 099;
            rddata_opt[2] <= 062;
            rddata_opt[3] <= 014;
          end
        0181: begin
            rddata_opt[0] <= 012;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 107;
          end
        0182: begin
            rddata_opt[0] <= 012;
            rddata_opt[1] <= 030;
            rddata_opt[2] <= 012;
            rddata_opt[3] <= 012;
          end
        0183: begin
            rddata_opt[0] <= 012;
            rddata_opt[1] <= 048;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0184: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 048;
            rddata_opt[2] <= 102;
            rddata_opt[3] <= 051;
          end
        0185: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 031;
            rddata_opt[3] <= 051;
          end
        0186: begin
            rddata_opt[0] <= 110;
            rddata_opt[1] <= 024;
            rddata_opt[2] <= 048;
            rddata_opt[3] <= 054;
          end
        0187: begin
            rddata_opt[0] <= 024;
            rddata_opt[1] <= 107;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 051;
          end
        0188: begin
            rddata_opt[0] <= 102;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 118;
            rddata_opt[3] <= 051;
          end
        0189: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 099;
          end
        0190: begin
            rddata_opt[0] <= 054;
            rddata_opt[1] <= 102;
            rddata_opt[2] <= 049;
            rddata_opt[3] <= 000;
          end
        0194: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 069;
            rddata_opt[3] <= 000;
          end
        0195: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 028;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0196: begin
            rddata_opt[0] <= 124;
            rddata_opt[1] <= 031;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0198: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 006;
            rddata_opt[3] <= 048;
          end
        0200: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0201: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0202: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 048;
            rddata_opt[2] <= 060;
            rddata_opt[3] <= 024;
          end
        0203: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 012;
          end
        0204: begin
            rddata_opt[0] <= 111;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 012;
            rddata_opt[3] <= 048;
          end
        0205: begin
            rddata_opt[0] <= 127;
            rddata_opt[1] <= 048;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 024;
          end
        0206: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 024;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0207: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 126;
            rddata_opt[2] <= 048;
            rddata_opt[3] <= 012;
          end
        0208: begin
            rddata_opt[0] <= 123;
            rddata_opt[1] <= 063;
            rddata_opt[2] <= 102;
            rddata_opt[3] <= 003;
          end
        0209: begin
            rddata_opt[0] <= 102;
            rddata_opt[1] <= 038;
            rddata_opt[2] <= 038;
            rddata_opt[3] <= 115;
          end
        0210: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 054;
          end
        0211: begin
            rddata_opt[0] <= 070;
            rddata_opt[1] <= 099;
            rddata_opt[2] <= 123;
            rddata_opt[3] <= 099;
          end
        0212: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 115;
            rddata_opt[2] <= 054;
            rddata_opt[3] <= 024;
          end
        0213: begin
            rddata_opt[0] <= 012;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 107;
          end
        0214: begin
            rddata_opt[0] <= 030;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 006;
            rddata_opt[3] <= 012;
          end
        0215: begin
            rddata_opt[0] <= 024;
            rddata_opt[1] <= 048;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0216: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 062;
            rddata_opt[2] <= 102;
            rddata_opt[3] <= 003;
          end
        0217: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 063;
            rddata_opt[2] <= 006;
            rddata_opt[3] <= 051;
          end
        0218: begin
            rddata_opt[0] <= 102;
            rddata_opt[1] <= 024;
            rddata_opt[2] <= 048;
            rddata_opt[3] <= 030;
          end
        0219: begin
            rddata_opt[0] <= 024;
            rddata_opt[1] <= 107;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 051;
          end
        0220: begin
            rddata_opt[0] <= 102;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 110;
            rddata_opt[3] <= 006;
          end
        0221: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 107;
          end
        0222: begin
            rddata_opt[0] <= 028;
            rddata_opt[1] <= 102;
            rddata_opt[2] <= 024;
            rddata_opt[3] <= 000;
          end
        0226: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 093;
            rddata_opt[3] <= 000;
          end
        0227: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 054;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0228: begin
            rddata_opt[0] <= 112;
            rddata_opt[1] <= 007;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0230: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 012;
            rddata_opt[3] <= 024;
          end
        0233: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 006;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0234: begin
            rddata_opt[0] <= 012;
            rddata_opt[1] <= 024;
            rddata_opt[2] <= 102;
            rddata_opt[3] <= 024;
          end
        0235: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 006;
          end
        0236: begin
            rddata_opt[0] <= 103;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 006;
            rddata_opt[3] <= 048;
          end
        0237: begin
            rddata_opt[0] <= 048;
            rddata_opt[1] <= 048;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 012;
          end
        0238: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 024;
            rddata_opt[2] <= 028;
            rddata_opt[3] <= 028;
          end
        0239: begin
            rddata_opt[0] <= 012;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 024;
            rddata_opt[3] <= 000;
          end
        0240: begin
            rddata_opt[0] <= 003;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 102;
            rddata_opt[3] <= 099;
          end
        0241: begin
            rddata_opt[0] <= 102;
            rddata_opt[1] <= 006;
            rddata_opt[2] <= 006;
            rddata_opt[3] <= 099;
          end
        0242: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 054;
          end
        0243: begin
            rddata_opt[0] <= 102;
            rddata_opt[1] <= 099;
            rddata_opt[2] <= 115;
            rddata_opt[3] <= 099;
          end
        0244: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 123;
            rddata_opt[2] <= 102;
            rddata_opt[3] <= 051;
          end
        0245: begin
            rddata_opt[0] <= 012;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 054;
          end
        0246: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 070;
            rddata_opt[3] <= 012;
          end
        0247: begin
            rddata_opt[0] <= 048;
            rddata_opt[1] <= 048;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0248: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 102;
            rddata_opt[3] <= 003;
          end
        0249: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 003;
            rddata_opt[2] <= 006;
            rddata_opt[3] <= 051;
          end
        0250: begin
            rddata_opt[0] <= 102;
            rddata_opt[1] <= 024;
            rddata_opt[2] <= 048;
            rddata_opt[3] <= 054;
          end
        0251: begin
            rddata_opt[0] <= 024;
            rddata_opt[1] <= 107;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 051;
          end
        0252: begin
            rddata_opt[0] <= 102;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 006;
            rddata_opt[3] <= 024;
          end
        0253: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 107;
          end
        0254: begin
            rddata_opt[0] <= 028;
            rddata_opt[1] <= 102;
            rddata_opt[2] <= 006;
            rddata_opt[3] <= 000;
          end
        0258: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 034;
            rddata_opt[3] <= 000;
          end
        0259: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 099;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0260: begin
            rddata_opt[0] <= 096;
            rddata_opt[1] <= 003;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0264: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0265: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0266: begin
            rddata_opt[0] <= 024;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0267: begin
            rddata_opt[0] <= 028;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 028;
            rddata_opt[3] <= 003;
          end
        0268: begin
            rddata_opt[0] <= 099;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 051;
          end
        0269: begin
            rddata_opt[0] <= 048;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 012;
          end
        0270: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 028;
            rddata_opt[3] <= 028;
          end
        0271: begin
            rddata_opt[0] <= 024;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 012;
            rddata_opt[3] <= 012;
          end
        0272: begin
            rddata_opt[0] <= 003;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 102;
            rddata_opt[3] <= 102;
          end
        0273: begin
            rddata_opt[0] <= 054;
            rddata_opt[1] <= 070;
            rddata_opt[2] <= 006;
            rddata_opt[3] <= 102;
          end
        0274: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 102;
          end
        0275: begin
            rddata_opt[0] <= 102;
            rddata_opt[1] <= 099;
            rddata_opt[2] <= 099;
            rddata_opt[3] <= 054;
          end
        0276: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 062;
            rddata_opt[2] <= 102;
            rddata_opt[3] <= 051;
          end
        0277: begin
            rddata_opt[0] <= 012;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 030;
            rddata_opt[3] <= 054;
          end
        0278: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 099;
            rddata_opt[3] <= 012;
          end
        0279: begin
            rddata_opt[0] <= 096;
            rddata_opt[1] <= 048;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0280: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 102;
            rddata_opt[3] <= 051;
          end
        0281: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 006;
            rddata_opt[3] <= 062;
          end
        0282: begin
            rddata_opt[0] <= 102;
            rddata_opt[1] <= 024;
            rddata_opt[2] <= 048;
            rddata_opt[3] <= 102;
          end
        0283: begin
            rddata_opt[0] <= 024;
            rddata_opt[1] <= 107;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 051;
          end
        0284: begin
            rddata_opt[0] <= 102;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 006;
            rddata_opt[3] <= 051;
          end
        0285: begin
            rddata_opt[0] <= 054;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 030;
            rddata_opt[3] <= 054;
          end
        0286: begin
            rddata_opt[0] <= 054;
            rddata_opt[1] <= 060;
            rddata_opt[2] <= 035;
            rddata_opt[3] <= 000;
          end
        0290: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 028;
            rddata_opt[3] <= 000;
          end
        0292: begin
            rddata_opt[0] <= 064;
            rddata_opt[1] <= 001;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0296: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 012;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0297: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 049;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0298: begin
            rddata_opt[0] <= 048;
            rddata_opt[1] <= 006;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0299: begin
            rddata_opt[0] <= 028;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 028;
            rddata_opt[3] <= 001;
          end
        0300: begin
            rddata_opt[0] <= 062;
            rddata_opt[1] <= 063;
            rddata_opt[2] <= 063;
            rddata_opt[3] <= 030;
          end
        0301: begin
            rddata_opt[0] <= 120;
            rddata_opt[1] <= 030;
            rddata_opt[2] <= 030;
            rddata_opt[3] <= 012;
          end
        0302: begin
            rddata_opt[0] <= 030;
            rddata_opt[1] <= 014;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 024;
          end
        0303: begin
            rddata_opt[0] <= 048;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 006;
            rddata_opt[3] <= 012;
          end
        0304: begin
            rddata_opt[0] <= 062;
            rddata_opt[1] <= 051;
            rddata_opt[2] <= 063;
            rddata_opt[3] <= 060;
          end
        0305: begin
            rddata_opt[0] <= 031;
            rddata_opt[1] <= 127;
            rddata_opt[2] <= 015;
            rddata_opt[3] <= 124;
          end
        0306: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 030;
            rddata_opt[2] <= 030;
            rddata_opt[3] <= 103;
          end
        0307: begin
            rddata_opt[0] <= 127;
            rddata_opt[1] <= 099;
            rddata_opt[2] <= 099;
            rddata_opt[3] <= 028;
          end
        0308: begin
            rddata_opt[0] <= 015;
            rddata_opt[1] <= 048;
            rddata_opt[2] <= 103;
            rddata_opt[3] <= 030;
          end
        0309: begin
            rddata_opt[0] <= 030;
            rddata_opt[1] <= 030;
            rddata_opt[2] <= 012;
            rddata_opt[3] <= 054;
          end
        0310: begin
            rddata_opt[0] <= 051;
            rddata_opt[1] <= 030;
            rddata_opt[2] <= 127;
            rddata_opt[3] <= 060;
          end
        0311: begin
            rddata_opt[0] <= 064;
            rddata_opt[1] <= 060;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0312: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 110;
            rddata_opt[2] <= 059;
            rddata_opt[3] <= 030;
          end
        0313: begin
            rddata_opt[0] <= 110;
            rddata_opt[1] <= 030;
            rddata_opt[2] <= 015;
            rddata_opt[3] <= 048;
          end
        0314: begin
            rddata_opt[0] <= 103;
            rddata_opt[1] <= 126;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 103;
          end
        0315: begin
            rddata_opt[0] <= 126;
            rddata_opt[1] <= 099;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 030;
          end
        0316: begin
            rddata_opt[0] <= 062;
            rddata_opt[1] <= 062;
            rddata_opt[2] <= 015;
            rddata_opt[3] <= 030;
          end
        0317: begin
            rddata_opt[0] <= 028;
            rddata_opt[1] <= 110;
            rddata_opt[2] <= 012;
            rddata_opt[3] <= 054;
          end
        0318: begin
            rddata_opt[0] <= 099;
            rddata_opt[1] <= 048;
            rddata_opt[2] <= 063;
            rddata_opt[3] <= 000;
          end
        0331: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0334: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 012;
          end
        0340: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 120;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0345: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 051;
          end
        0346: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 051;
            rddata_opt[3] <= 000;
          end
        0348: begin
            rddata_opt[0] <= 006;
            rddata_opt[1] <= 048;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0350: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 024;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0377: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 030;
          end
        0378: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 030;
            rddata_opt[3] <= 000;
          end
        0380: begin
            rddata_opt[0] <= 015;
            rddata_opt[1] <= 120;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        0382: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 015;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
        default: begin
            rddata_opt[0] <= 000;
            rddata_opt[1] <= 000;
            rddata_opt[2] <= 000;
            rddata_opt[3] <= 000;
          end
      endcase
    end
    if (rden_r)
      rddata <= rddata_opt[lsb_addr_r];
    end

endmodule
