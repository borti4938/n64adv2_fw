//////////////////////////////////////////////////////////////////////////////////
//
// This file is part of the N64 RGB/YPbPr DAC project.
//
// Copyright (C) 2015-2023 by Peter Bartmann <borti4938@gmail.com>
//
// N64 RGB/YPbPr DAC is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <http://www.gnu.org/licenses/>.
//
//////////////////////////////////////////////////////////////////////////////////
//
// Company:  Circuit-Board.de
// Engineer: borti4938
//
// Module Name:    gamma_table_v2
// Project Name:   N64 Advanced RGB/YPbPr DAC Mod
// Target Devices: universial
// Tool versions:  Altera Quartus Prime
// Description:    
//
// Features: ip independent implementation of gamma rom
//
// This file is auto generated by script/gamma2rom.m
//
//////////////////////////////////////////////////////////////////////////////////


module gamma_table_v2(
  VCLK,
  nRST,
  gamma_val,
  vdata_in,
  nbypass,
  vdata_out
);

`include "../../lib/n64adv_vparams.vh"

input                     VCLK;
input                     nRST;
input [              2:0] gamma_val;
input [color_width_i-1:0] vdata_in;
input                     nbypass;

output reg [color_width_o-1:0] vdata_out = {color_width_o{1'b0}};


reg [color_width_i+2:0] addr_r = {(color_width_i+3){1'b0}};
reg                  nbypass_r =  1'b0;

always @(posedge VCLK or negedge nRST)
  if (!nRST) begin
    vdata_out <= {(color_width_o){1'b0}};
       addr_r <= {(color_width_i+3){1'b0}};
    nbypass_r <=  1'b0;
  end else begin
    addr_r <= {gamma_val,vdata_in};
    nbypass_r <= nbypass;

    case (addr_r)
      0000: vdata_out <= 000;
      0001: vdata_out <= 007;
      0002: vdata_out <= 011;
      0003: vdata_out <= 015;
      0004: vdata_out <= 019;
      0005: vdata_out <= 023;
      0006: vdata_out <= 026;
      0007: vdata_out <= 029;
      0008: vdata_out <= 032;
      0009: vdata_out <= 035;
      0010: vdata_out <= 038;
      0011: vdata_out <= 041;
      0012: vdata_out <= 043;
      0013: vdata_out <= 046;
      0014: vdata_out <= 049;
      0015: vdata_out <= 051;
      0016: vdata_out <= 054;
      0017: vdata_out <= 056;
      0018: vdata_out <= 059;
      0019: vdata_out <= 061;
      0020: vdata_out <= 064;
      0021: vdata_out <= 066;
      0022: vdata_out <= 068;
      0023: vdata_out <= 071;
      0024: vdata_out <= 073;
      0025: vdata_out <= 075;
      0026: vdata_out <= 078;
      0027: vdata_out <= 080;
      0028: vdata_out <= 082;
      0029: vdata_out <= 084;
      0030: vdata_out <= 086;
      0031: vdata_out <= 089;
      0032: vdata_out <= 091;
      0033: vdata_out <= 093;
      0034: vdata_out <= 095;
      0035: vdata_out <= 097;
      0036: vdata_out <= 099;
      0037: vdata_out <= 101;
      0038: vdata_out <= 103;
      0039: vdata_out <= 105;
      0040: vdata_out <= 107;
      0041: vdata_out <= 109;
      0042: vdata_out <= 111;
      0043: vdata_out <= 113;
      0044: vdata_out <= 115;
      0045: vdata_out <= 117;
      0046: vdata_out <= 119;
      0047: vdata_out <= 121;
      0048: vdata_out <= 123;
      0049: vdata_out <= 125;
      0050: vdata_out <= 127;
      0051: vdata_out <= 129;
      0052: vdata_out <= 131;
      0053: vdata_out <= 132;
      0054: vdata_out <= 134;
      0055: vdata_out <= 136;
      0056: vdata_out <= 138;
      0057: vdata_out <= 140;
      0058: vdata_out <= 142;
      0059: vdata_out <= 143;
      0060: vdata_out <= 145;
      0061: vdata_out <= 147;
      0062: vdata_out <= 149;
      0063: vdata_out <= 151;
      0064: vdata_out <= 153;
      0065: vdata_out <= 154;
      0066: vdata_out <= 156;
      0067: vdata_out <= 158;
      0068: vdata_out <= 160;
      0069: vdata_out <= 161;
      0070: vdata_out <= 163;
      0071: vdata_out <= 165;
      0072: vdata_out <= 167;
      0073: vdata_out <= 168;
      0074: vdata_out <= 170;
      0075: vdata_out <= 172;
      0076: vdata_out <= 173;
      0077: vdata_out <= 175;
      0078: vdata_out <= 177;
      0079: vdata_out <= 179;
      0080: vdata_out <= 180;
      0081: vdata_out <= 182;
      0082: vdata_out <= 184;
      0083: vdata_out <= 185;
      0084: vdata_out <= 187;
      0085: vdata_out <= 189;
      0086: vdata_out <= 190;
      0087: vdata_out <= 192;
      0088: vdata_out <= 194;
      0089: vdata_out <= 195;
      0090: vdata_out <= 197;
      0091: vdata_out <= 199;
      0092: vdata_out <= 200;
      0093: vdata_out <= 202;
      0094: vdata_out <= 203;
      0095: vdata_out <= 205;
      0096: vdata_out <= 207;
      0097: vdata_out <= 208;
      0098: vdata_out <= 210;
      0099: vdata_out <= 212;
      0100: vdata_out <= 213;
      0101: vdata_out <= 215;
      0102: vdata_out <= 216;
      0103: vdata_out <= 218;
      0104: vdata_out <= 220;
      0105: vdata_out <= 221;
      0106: vdata_out <= 223;
      0107: vdata_out <= 224;
      0108: vdata_out <= 226;
      0109: vdata_out <= 227;
      0110: vdata_out <= 229;
      0111: vdata_out <= 231;
      0112: vdata_out <= 232;
      0113: vdata_out <= 234;
      0114: vdata_out <= 235;
      0115: vdata_out <= 237;
      0116: vdata_out <= 238;
      0117: vdata_out <= 240;
      0118: vdata_out <= 241;
      0119: vdata_out <= 243;
      0120: vdata_out <= 244;
      0121: vdata_out <= 246;
      0122: vdata_out <= 247;
      0123: vdata_out <= 249;
      0124: vdata_out <= 250;
      0125: vdata_out <= 252;
      0126: vdata_out <= 253;
      0127: vdata_out <= 255;
      0128: vdata_out <= 000;
      0129: vdata_out <= 005;
      0130: vdata_out <= 009;
      0131: vdata_out <= 013;
      0132: vdata_out <= 016;
      0133: vdata_out <= 019;
      0134: vdata_out <= 022;
      0135: vdata_out <= 025;
      0136: vdata_out <= 028;
      0137: vdata_out <= 031;
      0138: vdata_out <= 033;
      0139: vdata_out <= 036;
      0140: vdata_out <= 039;
      0141: vdata_out <= 041;
      0142: vdata_out <= 044;
      0143: vdata_out <= 046;
      0144: vdata_out <= 049;
      0145: vdata_out <= 051;
      0146: vdata_out <= 053;
      0147: vdata_out <= 056;
      0148: vdata_out <= 058;
      0149: vdata_out <= 060;
      0150: vdata_out <= 063;
      0151: vdata_out <= 065;
      0152: vdata_out <= 067;
      0153: vdata_out <= 069;
      0154: vdata_out <= 072;
      0155: vdata_out <= 074;
      0156: vdata_out <= 076;
      0157: vdata_out <= 078;
      0158: vdata_out <= 080;
      0159: vdata_out <= 083;
      0160: vdata_out <= 085;
      0161: vdata_out <= 087;
      0162: vdata_out <= 089;
      0163: vdata_out <= 091;
      0164: vdata_out <= 093;
      0165: vdata_out <= 095;
      0166: vdata_out <= 097;
      0167: vdata_out <= 099;
      0168: vdata_out <= 101;
      0169: vdata_out <= 103;
      0170: vdata_out <= 105;
      0171: vdata_out <= 107;
      0172: vdata_out <= 109;
      0173: vdata_out <= 111;
      0174: vdata_out <= 113;
      0175: vdata_out <= 115;
      0176: vdata_out <= 117;
      0177: vdata_out <= 119;
      0178: vdata_out <= 121;
      0179: vdata_out <= 123;
      0180: vdata_out <= 125;
      0181: vdata_out <= 127;
      0182: vdata_out <= 129;
      0183: vdata_out <= 131;
      0184: vdata_out <= 132;
      0185: vdata_out <= 134;
      0186: vdata_out <= 136;
      0187: vdata_out <= 138;
      0188: vdata_out <= 140;
      0189: vdata_out <= 142;
      0190: vdata_out <= 144;
      0191: vdata_out <= 146;
      0192: vdata_out <= 147;
      0193: vdata_out <= 149;
      0194: vdata_out <= 151;
      0195: vdata_out <= 153;
      0196: vdata_out <= 155;
      0197: vdata_out <= 157;
      0198: vdata_out <= 158;
      0199: vdata_out <= 160;
      0200: vdata_out <= 162;
      0201: vdata_out <= 164;
      0202: vdata_out <= 166;
      0203: vdata_out <= 167;
      0204: vdata_out <= 169;
      0205: vdata_out <= 171;
      0206: vdata_out <= 173;
      0207: vdata_out <= 174;
      0208: vdata_out <= 176;
      0209: vdata_out <= 178;
      0210: vdata_out <= 180;
      0211: vdata_out <= 181;
      0212: vdata_out <= 183;
      0213: vdata_out <= 185;
      0214: vdata_out <= 187;
      0215: vdata_out <= 188;
      0216: vdata_out <= 190;
      0217: vdata_out <= 192;
      0218: vdata_out <= 194;
      0219: vdata_out <= 195;
      0220: vdata_out <= 197;
      0221: vdata_out <= 199;
      0222: vdata_out <= 200;
      0223: vdata_out <= 202;
      0224: vdata_out <= 204;
      0225: vdata_out <= 206;
      0226: vdata_out <= 207;
      0227: vdata_out <= 209;
      0228: vdata_out <= 211;
      0229: vdata_out <= 212;
      0230: vdata_out <= 214;
      0231: vdata_out <= 216;
      0232: vdata_out <= 217;
      0233: vdata_out <= 219;
      0234: vdata_out <= 221;
      0235: vdata_out <= 222;
      0236: vdata_out <= 224;
      0237: vdata_out <= 226;
      0238: vdata_out <= 227;
      0239: vdata_out <= 229;
      0240: vdata_out <= 231;
      0241: vdata_out <= 232;
      0242: vdata_out <= 234;
      0243: vdata_out <= 236;
      0244: vdata_out <= 237;
      0245: vdata_out <= 239;
      0246: vdata_out <= 240;
      0247: vdata_out <= 242;
      0248: vdata_out <= 244;
      0249: vdata_out <= 245;
      0250: vdata_out <= 247;
      0251: vdata_out <= 249;
      0252: vdata_out <= 250;
      0253: vdata_out <= 252;
      0254: vdata_out <= 253;
      0255: vdata_out <= 255;
      0256: vdata_out <= 000;
      0257: vdata_out <= 004;
      0258: vdata_out <= 007;
      0259: vdata_out <= 011;
      0260: vdata_out <= 013;
      0261: vdata_out <= 016;
      0262: vdata_out <= 019;
      0263: vdata_out <= 022;
      0264: vdata_out <= 024;
      0265: vdata_out <= 027;
      0266: vdata_out <= 029;
      0267: vdata_out <= 032;
      0268: vdata_out <= 034;
      0269: vdata_out <= 037;
      0270: vdata_out <= 039;
      0271: vdata_out <= 041;
      0272: vdata_out <= 044;
      0273: vdata_out <= 046;
      0274: vdata_out <= 048;
      0275: vdata_out <= 051;
      0276: vdata_out <= 053;
      0277: vdata_out <= 055;
      0278: vdata_out <= 057;
      0279: vdata_out <= 060;
      0280: vdata_out <= 062;
      0281: vdata_out <= 064;
      0282: vdata_out <= 066;
      0283: vdata_out <= 068;
      0284: vdata_out <= 071;
      0285: vdata_out <= 073;
      0286: vdata_out <= 075;
      0287: vdata_out <= 077;
      0288: vdata_out <= 079;
      0289: vdata_out <= 081;
      0290: vdata_out <= 083;
      0291: vdata_out <= 085;
      0292: vdata_out <= 087;
      0293: vdata_out <= 089;
      0294: vdata_out <= 091;
      0295: vdata_out <= 093;
      0296: vdata_out <= 096;
      0297: vdata_out <= 098;
      0298: vdata_out <= 100;
      0299: vdata_out <= 102;
      0300: vdata_out <= 104;
      0301: vdata_out <= 106;
      0302: vdata_out <= 108;
      0303: vdata_out <= 110;
      0304: vdata_out <= 112;
      0305: vdata_out <= 113;
      0306: vdata_out <= 115;
      0307: vdata_out <= 117;
      0308: vdata_out <= 119;
      0309: vdata_out <= 121;
      0310: vdata_out <= 123;
      0311: vdata_out <= 125;
      0312: vdata_out <= 127;
      0313: vdata_out <= 129;
      0314: vdata_out <= 131;
      0315: vdata_out <= 133;
      0316: vdata_out <= 135;
      0317: vdata_out <= 137;
      0318: vdata_out <= 139;
      0319: vdata_out <= 141;
      0320: vdata_out <= 142;
      0321: vdata_out <= 144;
      0322: vdata_out <= 146;
      0323: vdata_out <= 148;
      0324: vdata_out <= 150;
      0325: vdata_out <= 152;
      0326: vdata_out <= 154;
      0327: vdata_out <= 156;
      0328: vdata_out <= 157;
      0329: vdata_out <= 159;
      0330: vdata_out <= 161;
      0331: vdata_out <= 163;
      0332: vdata_out <= 165;
      0333: vdata_out <= 167;
      0334: vdata_out <= 168;
      0335: vdata_out <= 170;
      0336: vdata_out <= 172;
      0337: vdata_out <= 174;
      0338: vdata_out <= 176;
      0339: vdata_out <= 178;
      0340: vdata_out <= 179;
      0341: vdata_out <= 181;
      0342: vdata_out <= 183;
      0343: vdata_out <= 185;
      0344: vdata_out <= 187;
      0345: vdata_out <= 188;
      0346: vdata_out <= 190;
      0347: vdata_out <= 192;
      0348: vdata_out <= 194;
      0349: vdata_out <= 196;
      0350: vdata_out <= 197;
      0351: vdata_out <= 199;
      0352: vdata_out <= 201;
      0353: vdata_out <= 203;
      0354: vdata_out <= 205;
      0355: vdata_out <= 206;
      0356: vdata_out <= 208;
      0357: vdata_out <= 210;
      0358: vdata_out <= 212;
      0359: vdata_out <= 213;
      0360: vdata_out <= 215;
      0361: vdata_out <= 217;
      0362: vdata_out <= 219;
      0363: vdata_out <= 220;
      0364: vdata_out <= 222;
      0365: vdata_out <= 224;
      0366: vdata_out <= 226;
      0367: vdata_out <= 227;
      0368: vdata_out <= 229;
      0369: vdata_out <= 231;
      0370: vdata_out <= 233;
      0371: vdata_out <= 234;
      0372: vdata_out <= 236;
      0373: vdata_out <= 238;
      0374: vdata_out <= 240;
      0375: vdata_out <= 241;
      0376: vdata_out <= 243;
      0377: vdata_out <= 245;
      0378: vdata_out <= 246;
      0379: vdata_out <= 248;
      0380: vdata_out <= 250;
      0381: vdata_out <= 252;
      0382: vdata_out <= 253;
      0383: vdata_out <= 255;
      0384: vdata_out <= 000;
      0385: vdata_out <= 003;
      0386: vdata_out <= 006;
      0387: vdata_out <= 009;
      0388: vdata_out <= 011;
      0389: vdata_out <= 014;
      0390: vdata_out <= 016;
      0391: vdata_out <= 019;
      0392: vdata_out <= 021;
      0393: vdata_out <= 024;
      0394: vdata_out <= 026;
      0395: vdata_out <= 028;
      0396: vdata_out <= 031;
      0397: vdata_out <= 033;
      0398: vdata_out <= 035;
      0399: vdata_out <= 037;
      0400: vdata_out <= 040;
      0401: vdata_out <= 042;
      0402: vdata_out <= 044;
      0403: vdata_out <= 046;
      0404: vdata_out <= 048;
      0405: vdata_out <= 050;
      0406: vdata_out <= 053;
      0407: vdata_out <= 055;
      0408: vdata_out <= 057;
      0409: vdata_out <= 059;
      0410: vdata_out <= 061;
      0411: vdata_out <= 063;
      0412: vdata_out <= 065;
      0413: vdata_out <= 067;
      0414: vdata_out <= 070;
      0415: vdata_out <= 072;
      0416: vdata_out <= 074;
      0417: vdata_out <= 076;
      0418: vdata_out <= 078;
      0419: vdata_out <= 080;
      0420: vdata_out <= 082;
      0421: vdata_out <= 084;
      0422: vdata_out <= 086;
      0423: vdata_out <= 088;
      0424: vdata_out <= 090;
      0425: vdata_out <= 092;
      0426: vdata_out <= 094;
      0427: vdata_out <= 096;
      0428: vdata_out <= 098;
      0429: vdata_out <= 100;
      0430: vdata_out <= 102;
      0431: vdata_out <= 104;
      0432: vdata_out <= 106;
      0433: vdata_out <= 108;
      0434: vdata_out <= 110;
      0435: vdata_out <= 112;
      0436: vdata_out <= 114;
      0437: vdata_out <= 116;
      0438: vdata_out <= 118;
      0439: vdata_out <= 120;
      0440: vdata_out <= 122;
      0441: vdata_out <= 124;
      0442: vdata_out <= 126;
      0443: vdata_out <= 128;
      0444: vdata_out <= 130;
      0445: vdata_out <= 132;
      0446: vdata_out <= 134;
      0447: vdata_out <= 136;
      0448: vdata_out <= 138;
      0449: vdata_out <= 140;
      0450: vdata_out <= 141;
      0451: vdata_out <= 143;
      0452: vdata_out <= 145;
      0453: vdata_out <= 147;
      0454: vdata_out <= 149;
      0455: vdata_out <= 151;
      0456: vdata_out <= 153;
      0457: vdata_out <= 155;
      0458: vdata_out <= 157;
      0459: vdata_out <= 159;
      0460: vdata_out <= 161;
      0461: vdata_out <= 163;
      0462: vdata_out <= 164;
      0463: vdata_out <= 166;
      0464: vdata_out <= 168;
      0465: vdata_out <= 170;
      0466: vdata_out <= 172;
      0467: vdata_out <= 174;
      0468: vdata_out <= 176;
      0469: vdata_out <= 178;
      0470: vdata_out <= 180;
      0471: vdata_out <= 181;
      0472: vdata_out <= 183;
      0473: vdata_out <= 185;
      0474: vdata_out <= 187;
      0475: vdata_out <= 189;
      0476: vdata_out <= 191;
      0477: vdata_out <= 193;
      0478: vdata_out <= 195;
      0479: vdata_out <= 196;
      0480: vdata_out <= 198;
      0481: vdata_out <= 200;
      0482: vdata_out <= 202;
      0483: vdata_out <= 204;
      0484: vdata_out <= 206;
      0485: vdata_out <= 207;
      0486: vdata_out <= 209;
      0487: vdata_out <= 211;
      0488: vdata_out <= 213;
      0489: vdata_out <= 215;
      0490: vdata_out <= 217;
      0491: vdata_out <= 219;
      0492: vdata_out <= 220;
      0493: vdata_out <= 222;
      0494: vdata_out <= 224;
      0495: vdata_out <= 226;
      0496: vdata_out <= 228;
      0497: vdata_out <= 230;
      0498: vdata_out <= 231;
      0499: vdata_out <= 233;
      0500: vdata_out <= 235;
      0501: vdata_out <= 237;
      0502: vdata_out <= 239;
      0503: vdata_out <= 240;
      0504: vdata_out <= 242;
      0505: vdata_out <= 244;
      0506: vdata_out <= 246;
      0507: vdata_out <= 248;
      0508: vdata_out <= 250;
      0509: vdata_out <= 251;
      0510: vdata_out <= 253;
      0511: vdata_out <= 255;
      0512: vdata_out <= 000;
      0513: vdata_out <= 003;
      0514: vdata_out <= 005;
      0515: vdata_out <= 007;
      0516: vdata_out <= 010;
      0517: vdata_out <= 012;
      0518: vdata_out <= 014;
      0519: vdata_out <= 016;
      0520: vdata_out <= 018;
      0521: vdata_out <= 021;
      0522: vdata_out <= 023;
      0523: vdata_out <= 025;
      0524: vdata_out <= 027;
      0525: vdata_out <= 029;
      0526: vdata_out <= 031;
      0527: vdata_out <= 034;
      0528: vdata_out <= 036;
      0529: vdata_out <= 038;
      0530: vdata_out <= 040;
      0531: vdata_out <= 042;
      0532: vdata_out <= 044;
      0533: vdata_out <= 046;
      0534: vdata_out <= 048;
      0535: vdata_out <= 050;
      0536: vdata_out <= 052;
      0537: vdata_out <= 054;
      0538: vdata_out <= 057;
      0539: vdata_out <= 059;
      0540: vdata_out <= 061;
      0541: vdata_out <= 063;
      0542: vdata_out <= 065;
      0543: vdata_out <= 067;
      0544: vdata_out <= 069;
      0545: vdata_out <= 071;
      0546: vdata_out <= 073;
      0547: vdata_out <= 075;
      0548: vdata_out <= 077;
      0549: vdata_out <= 079;
      0550: vdata_out <= 081;
      0551: vdata_out <= 083;
      0552: vdata_out <= 085;
      0553: vdata_out <= 087;
      0554: vdata_out <= 089;
      0555: vdata_out <= 091;
      0556: vdata_out <= 093;
      0557: vdata_out <= 095;
      0558: vdata_out <= 097;
      0559: vdata_out <= 099;
      0560: vdata_out <= 101;
      0561: vdata_out <= 103;
      0562: vdata_out <= 105;
      0563: vdata_out <= 107;
      0564: vdata_out <= 109;
      0565: vdata_out <= 111;
      0566: vdata_out <= 113;
      0567: vdata_out <= 115;
      0568: vdata_out <= 117;
      0569: vdata_out <= 119;
      0570: vdata_out <= 121;
      0571: vdata_out <= 123;
      0572: vdata_out <= 125;
      0573: vdata_out <= 127;
      0574: vdata_out <= 129;
      0575: vdata_out <= 131;
      0576: vdata_out <= 133;
      0577: vdata_out <= 135;
      0578: vdata_out <= 137;
      0579: vdata_out <= 139;
      0580: vdata_out <= 141;
      0581: vdata_out <= 143;
      0582: vdata_out <= 145;
      0583: vdata_out <= 147;
      0584: vdata_out <= 149;
      0585: vdata_out <= 151;
      0586: vdata_out <= 153;
      0587: vdata_out <= 155;
      0588: vdata_out <= 157;
      0589: vdata_out <= 159;
      0590: vdata_out <= 160;
      0591: vdata_out <= 162;
      0592: vdata_out <= 164;
      0593: vdata_out <= 166;
      0594: vdata_out <= 168;
      0595: vdata_out <= 170;
      0596: vdata_out <= 172;
      0597: vdata_out <= 174;
      0598: vdata_out <= 176;
      0599: vdata_out <= 178;
      0600: vdata_out <= 180;
      0601: vdata_out <= 182;
      0602: vdata_out <= 184;
      0603: vdata_out <= 186;
      0604: vdata_out <= 188;
      0605: vdata_out <= 190;
      0606: vdata_out <= 192;
      0607: vdata_out <= 194;
      0608: vdata_out <= 195;
      0609: vdata_out <= 197;
      0610: vdata_out <= 199;
      0611: vdata_out <= 201;
      0612: vdata_out <= 203;
      0613: vdata_out <= 205;
      0614: vdata_out <= 207;
      0615: vdata_out <= 209;
      0616: vdata_out <= 211;
      0617: vdata_out <= 213;
      0618: vdata_out <= 215;
      0619: vdata_out <= 217;
      0620: vdata_out <= 219;
      0621: vdata_out <= 221;
      0622: vdata_out <= 222;
      0623: vdata_out <= 224;
      0624: vdata_out <= 226;
      0625: vdata_out <= 228;
      0626: vdata_out <= 230;
      0627: vdata_out <= 232;
      0628: vdata_out <= 234;
      0629: vdata_out <= 236;
      0630: vdata_out <= 238;
      0631: vdata_out <= 240;
      0632: vdata_out <= 242;
      0633: vdata_out <= 244;
      0634: vdata_out <= 245;
      0635: vdata_out <= 247;
      0636: vdata_out <= 249;
      0637: vdata_out <= 251;
      0638: vdata_out <= 253;
      0639: vdata_out <= 255;
      0640: vdata_out <= 000;
      0641: vdata_out <= 002;
      0642: vdata_out <= 003;
      0643: vdata_out <= 005;
      0644: vdata_out <= 007;
      0645: vdata_out <= 009;
      0646: vdata_out <= 010;
      0647: vdata_out <= 012;
      0648: vdata_out <= 014;
      0649: vdata_out <= 016;
      0650: vdata_out <= 018;
      0651: vdata_out <= 020;
      0652: vdata_out <= 021;
      0653: vdata_out <= 023;
      0654: vdata_out <= 025;
      0655: vdata_out <= 027;
      0656: vdata_out <= 029;
      0657: vdata_out <= 031;
      0658: vdata_out <= 033;
      0659: vdata_out <= 035;
      0660: vdata_out <= 037;
      0661: vdata_out <= 039;
      0662: vdata_out <= 040;
      0663: vdata_out <= 042;
      0664: vdata_out <= 044;
      0665: vdata_out <= 046;
      0666: vdata_out <= 048;
      0667: vdata_out <= 050;
      0668: vdata_out <= 052;
      0669: vdata_out <= 054;
      0670: vdata_out <= 056;
      0671: vdata_out <= 058;
      0672: vdata_out <= 060;
      0673: vdata_out <= 062;
      0674: vdata_out <= 064;
      0675: vdata_out <= 066;
      0676: vdata_out <= 068;
      0677: vdata_out <= 070;
      0678: vdata_out <= 072;
      0679: vdata_out <= 074;
      0680: vdata_out <= 076;
      0681: vdata_out <= 078;
      0682: vdata_out <= 080;
      0683: vdata_out <= 082;
      0684: vdata_out <= 084;
      0685: vdata_out <= 086;
      0686: vdata_out <= 088;
      0687: vdata_out <= 090;
      0688: vdata_out <= 092;
      0689: vdata_out <= 094;
      0690: vdata_out <= 096;
      0691: vdata_out <= 098;
      0692: vdata_out <= 100;
      0693: vdata_out <= 102;
      0694: vdata_out <= 104;
      0695: vdata_out <= 106;
      0696: vdata_out <= 108;
      0697: vdata_out <= 110;
      0698: vdata_out <= 112;
      0699: vdata_out <= 114;
      0700: vdata_out <= 116;
      0701: vdata_out <= 118;
      0702: vdata_out <= 120;
      0703: vdata_out <= 122;
      0704: vdata_out <= 124;
      0705: vdata_out <= 126;
      0706: vdata_out <= 128;
      0707: vdata_out <= 130;
      0708: vdata_out <= 132;
      0709: vdata_out <= 134;
      0710: vdata_out <= 136;
      0711: vdata_out <= 138;
      0712: vdata_out <= 141;
      0713: vdata_out <= 143;
      0714: vdata_out <= 145;
      0715: vdata_out <= 147;
      0716: vdata_out <= 149;
      0717: vdata_out <= 151;
      0718: vdata_out <= 153;
      0719: vdata_out <= 155;
      0720: vdata_out <= 157;
      0721: vdata_out <= 159;
      0722: vdata_out <= 161;
      0723: vdata_out <= 163;
      0724: vdata_out <= 165;
      0725: vdata_out <= 167;
      0726: vdata_out <= 169;
      0727: vdata_out <= 171;
      0728: vdata_out <= 173;
      0729: vdata_out <= 176;
      0730: vdata_out <= 178;
      0731: vdata_out <= 180;
      0732: vdata_out <= 182;
      0733: vdata_out <= 184;
      0734: vdata_out <= 186;
      0735: vdata_out <= 188;
      0736: vdata_out <= 190;
      0737: vdata_out <= 192;
      0738: vdata_out <= 194;
      0739: vdata_out <= 196;
      0740: vdata_out <= 198;
      0741: vdata_out <= 200;
      0742: vdata_out <= 203;
      0743: vdata_out <= 205;
      0744: vdata_out <= 207;
      0745: vdata_out <= 209;
      0746: vdata_out <= 211;
      0747: vdata_out <= 213;
      0748: vdata_out <= 215;
      0749: vdata_out <= 217;
      0750: vdata_out <= 219;
      0751: vdata_out <= 221;
      0752: vdata_out <= 223;
      0753: vdata_out <= 226;
      0754: vdata_out <= 228;
      0755: vdata_out <= 230;
      0756: vdata_out <= 232;
      0757: vdata_out <= 234;
      0758: vdata_out <= 236;
      0759: vdata_out <= 238;
      0760: vdata_out <= 240;
      0761: vdata_out <= 242;
      0762: vdata_out <= 244;
      0763: vdata_out <= 247;
      0764: vdata_out <= 249;
      0765: vdata_out <= 251;
      0766: vdata_out <= 253;
      0767: vdata_out <= 255;
      0768: vdata_out <= 000;
      0769: vdata_out <= 001;
      0770: vdata_out <= 003;
      0771: vdata_out <= 004;
      0772: vdata_out <= 006;
      0773: vdata_out <= 007;
      0774: vdata_out <= 009;
      0775: vdata_out <= 011;
      0776: vdata_out <= 012;
      0777: vdata_out <= 014;
      0778: vdata_out <= 016;
      0779: vdata_out <= 017;
      0780: vdata_out <= 019;
      0781: vdata_out <= 021;
      0782: vdata_out <= 023;
      0783: vdata_out <= 024;
      0784: vdata_out <= 026;
      0785: vdata_out <= 028;
      0786: vdata_out <= 030;
      0787: vdata_out <= 032;
      0788: vdata_out <= 033;
      0789: vdata_out <= 035;
      0790: vdata_out <= 037;
      0791: vdata_out <= 039;
      0792: vdata_out <= 041;
      0793: vdata_out <= 043;
      0794: vdata_out <= 045;
      0795: vdata_out <= 046;
      0796: vdata_out <= 048;
      0797: vdata_out <= 050;
      0798: vdata_out <= 052;
      0799: vdata_out <= 054;
      0800: vdata_out <= 056;
      0801: vdata_out <= 058;
      0802: vdata_out <= 060;
      0803: vdata_out <= 062;
      0804: vdata_out <= 064;
      0805: vdata_out <= 066;
      0806: vdata_out <= 068;
      0807: vdata_out <= 070;
      0808: vdata_out <= 072;
      0809: vdata_out <= 074;
      0810: vdata_out <= 075;
      0811: vdata_out <= 077;
      0812: vdata_out <= 079;
      0813: vdata_out <= 081;
      0814: vdata_out <= 083;
      0815: vdata_out <= 085;
      0816: vdata_out <= 087;
      0817: vdata_out <= 089;
      0818: vdata_out <= 091;
      0819: vdata_out <= 093;
      0820: vdata_out <= 095;
      0821: vdata_out <= 098;
      0822: vdata_out <= 100;
      0823: vdata_out <= 102;
      0824: vdata_out <= 104;
      0825: vdata_out <= 106;
      0826: vdata_out <= 108;
      0827: vdata_out <= 110;
      0828: vdata_out <= 112;
      0829: vdata_out <= 114;
      0830: vdata_out <= 116;
      0831: vdata_out <= 118;
      0832: vdata_out <= 120;
      0833: vdata_out <= 122;
      0834: vdata_out <= 124;
      0835: vdata_out <= 126;
      0836: vdata_out <= 128;
      0837: vdata_out <= 130;
      0838: vdata_out <= 132;
      0839: vdata_out <= 135;
      0840: vdata_out <= 137;
      0841: vdata_out <= 139;
      0842: vdata_out <= 141;
      0843: vdata_out <= 143;
      0844: vdata_out <= 145;
      0845: vdata_out <= 147;
      0846: vdata_out <= 149;
      0847: vdata_out <= 151;
      0848: vdata_out <= 153;
      0849: vdata_out <= 155;
      0850: vdata_out <= 158;
      0851: vdata_out <= 160;
      0852: vdata_out <= 162;
      0853: vdata_out <= 164;
      0854: vdata_out <= 166;
      0855: vdata_out <= 168;
      0856: vdata_out <= 170;
      0857: vdata_out <= 172;
      0858: vdata_out <= 175;
      0859: vdata_out <= 177;
      0860: vdata_out <= 179;
      0861: vdata_out <= 181;
      0862: vdata_out <= 183;
      0863: vdata_out <= 185;
      0864: vdata_out <= 187;
      0865: vdata_out <= 190;
      0866: vdata_out <= 192;
      0867: vdata_out <= 194;
      0868: vdata_out <= 196;
      0869: vdata_out <= 198;
      0870: vdata_out <= 200;
      0871: vdata_out <= 203;
      0872: vdata_out <= 205;
      0873: vdata_out <= 207;
      0874: vdata_out <= 209;
      0875: vdata_out <= 211;
      0876: vdata_out <= 213;
      0877: vdata_out <= 216;
      0878: vdata_out <= 218;
      0879: vdata_out <= 220;
      0880: vdata_out <= 222;
      0881: vdata_out <= 224;
      0882: vdata_out <= 226;
      0883: vdata_out <= 229;
      0884: vdata_out <= 231;
      0885: vdata_out <= 233;
      0886: vdata_out <= 235;
      0887: vdata_out <= 237;
      0888: vdata_out <= 240;
      0889: vdata_out <= 242;
      0890: vdata_out <= 244;
      0891: vdata_out <= 246;
      0892: vdata_out <= 248;
      0893: vdata_out <= 251;
      0894: vdata_out <= 253;
      0895: vdata_out <= 255;
      0896: vdata_out <= 000;
      0897: vdata_out <= 001;
      0898: vdata_out <= 002;
      0899: vdata_out <= 003;
      0900: vdata_out <= 005;
      0901: vdata_out <= 006;
      0902: vdata_out <= 008;
      0903: vdata_out <= 009;
      0904: vdata_out <= 011;
      0905: vdata_out <= 012;
      0906: vdata_out <= 014;
      0907: vdata_out <= 015;
      0908: vdata_out <= 017;
      0909: vdata_out <= 019;
      0910: vdata_out <= 020;
      0911: vdata_out <= 022;
      0912: vdata_out <= 024;
      0913: vdata_out <= 025;
      0914: vdata_out <= 027;
      0915: vdata_out <= 029;
      0916: vdata_out <= 030;
      0917: vdata_out <= 032;
      0918: vdata_out <= 034;
      0919: vdata_out <= 036;
      0920: vdata_out <= 038;
      0921: vdata_out <= 039;
      0922: vdata_out <= 041;
      0923: vdata_out <= 043;
      0924: vdata_out <= 045;
      0925: vdata_out <= 047;
      0926: vdata_out <= 049;
      0927: vdata_out <= 050;
      0928: vdata_out <= 052;
      0929: vdata_out <= 054;
      0930: vdata_out <= 056;
      0931: vdata_out <= 058;
      0932: vdata_out <= 060;
      0933: vdata_out <= 062;
      0934: vdata_out <= 064;
      0935: vdata_out <= 066;
      0936: vdata_out <= 068;
      0937: vdata_out <= 069;
      0938: vdata_out <= 071;
      0939: vdata_out <= 073;
      0940: vdata_out <= 075;
      0941: vdata_out <= 077;
      0942: vdata_out <= 079;
      0943: vdata_out <= 081;
      0944: vdata_out <= 083;
      0945: vdata_out <= 085;
      0946: vdata_out <= 087;
      0947: vdata_out <= 089;
      0948: vdata_out <= 091;
      0949: vdata_out <= 093;
      0950: vdata_out <= 095;
      0951: vdata_out <= 097;
      0952: vdata_out <= 099;
      0953: vdata_out <= 101;
      0954: vdata_out <= 104;
      0955: vdata_out <= 106;
      0956: vdata_out <= 108;
      0957: vdata_out <= 110;
      0958: vdata_out <= 112;
      0959: vdata_out <= 114;
      0960: vdata_out <= 116;
      0961: vdata_out <= 118;
      0962: vdata_out <= 120;
      0963: vdata_out <= 122;
      0964: vdata_out <= 124;
      0965: vdata_out <= 126;
      0966: vdata_out <= 129;
      0967: vdata_out <= 131;
      0968: vdata_out <= 133;
      0969: vdata_out <= 135;
      0970: vdata_out <= 137;
      0971: vdata_out <= 139;
      0972: vdata_out <= 141;
      0973: vdata_out <= 143;
      0974: vdata_out <= 146;
      0975: vdata_out <= 148;
      0976: vdata_out <= 150;
      0977: vdata_out <= 152;
      0978: vdata_out <= 154;
      0979: vdata_out <= 156;
      0980: vdata_out <= 159;
      0981: vdata_out <= 161;
      0982: vdata_out <= 163;
      0983: vdata_out <= 165;
      0984: vdata_out <= 167;
      0985: vdata_out <= 169;
      0986: vdata_out <= 172;
      0987: vdata_out <= 174;
      0988: vdata_out <= 176;
      0989: vdata_out <= 178;
      0990: vdata_out <= 180;
      0991: vdata_out <= 183;
      0992: vdata_out <= 185;
      0993: vdata_out <= 187;
      0994: vdata_out <= 189;
      0995: vdata_out <= 191;
      0996: vdata_out <= 194;
      0997: vdata_out <= 196;
      0998: vdata_out <= 198;
      0999: vdata_out <= 200;
      1000: vdata_out <= 203;
      1001: vdata_out <= 205;
      1002: vdata_out <= 207;
      1003: vdata_out <= 209;
      1004: vdata_out <= 212;
      1005: vdata_out <= 214;
      1006: vdata_out <= 216;
      1007: vdata_out <= 218;
      1008: vdata_out <= 221;
      1009: vdata_out <= 223;
      1010: vdata_out <= 225;
      1011: vdata_out <= 227;
      1012: vdata_out <= 230;
      1013: vdata_out <= 232;
      1014: vdata_out <= 234;
      1015: vdata_out <= 237;
      1016: vdata_out <= 239;
      1017: vdata_out <= 241;
      1018: vdata_out <= 243;
      1019: vdata_out <= 246;
      1020: vdata_out <= 248;
      1021: vdata_out <= 250;
      1022: vdata_out <= 253;
      1023: vdata_out <= 255;
    endcase

    if (!nbypass_r)
      vdata_out <= {addr_r[color_width_i-1:0],{1{vdata_in[color_width_i-1]}}};
  end

endmodule
